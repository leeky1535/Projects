module songdata(input logic clk,
					 input logic [12:0] addr,
					 output logic [3:0] data);
					 
reg [3:0] notes [0:255];

initial begin

		notes[0] = 4'b0000;  //measure 0
		notes[1] = 4'b0000;
		notes[2] = 4'b0000;
		notes[3] = 4'b0000;
		notes[4] = 4'b0000;  //measure 1
		notes[5] = 4'b1000;
		notes[6] = 4'b0000;
		notes[7] = 4'b0001;
		notes[8] = 4'b0000;  //measure 2
		notes[9] = 4'b1000;
		notes[10] = 4'b0000;
		notes[11] = 4'b0010;
		notes[12] = 4'b1000;  //measure 3
		notes[13] = 4'b0100;
		notes[14] = 4'b0000;
		notes[15] = 4'b0001;
		notes[16] = 4'b0000;  //measure 4
		notes[17] = 4'b1000;
		notes[18] = 4'b0000;
		notes[19] = 4'b0010;
		notes[20] = 4'b0000;  //measure 5
		notes[21] = 4'b1000;
		notes[22] = 4'b0000;
		notes[23] = 4'b0100;
		notes[24] = 4'b0000;  //measure 6
		notes[25] = 4'b0010;
		notes[26] = 4'b0000;
		notes[27] = 4'b0100;
		notes[28] = 4'b1000;  //measure 7
		notes[29] = 4'b0001;
		notes[30] = 4'b0000;
		notes[31] = 4'b0001;
		notes[32] = 4'b0000;  //measure 8
		notes[33] = 4'b0000;
		notes[34] = 4'b0000;
		notes[35] = 4'b0000;
		notes[36] = 4'b0000;  //measure 9
		notes[37] = 4'b1000;
		notes[38] = 4'b0001;
		notes[39] = 4'b1000;
		notes[40] = 4'b0010;  //measure 10
		notes[41] = 4'b0100;
		notes[42] = 4'b0001;
		notes[43] = 4'b0100;
		notes[44] = 4'b0100;  //measure 11
		notes[45] = 4'b0001;
		notes[46] = 4'b0100;
		notes[47] = 4'b0010;
		notes[48] = 4'b1000;  //measure 12
		notes[49] = 4'b0001;
		notes[50] = 4'b0000;
		notes[51] = 4'b0000;
		notes[52] = 4'b0000;  //measure 13
		notes[53] = 4'b0000;
		notes[54] = 4'b0000;
		notes[55] = 4'b0000;
		notes[56] = 4'b0001;  //measure 14
		notes[57] = 4'b0001;
		notes[58] = 4'b1000;
		notes[59] = 4'b0010;
		notes[60] = 4'b0100;  //measure 15
		notes[61] = 4'b0010;
		notes[62] = 4'b0000;
		notes[63] = 4'b0000;
		notes[64] = 4'b0010;  //measure 16
		notes[65] = 4'b0100;
		notes[66] = 4'b0001;
		notes[67] = 4'b0010;
		notes[68] = 4'b1000;  //measure 17
		notes[69] = 4'b0001;
		notes[70] = 4'b0000;
		notes[71] = 4'b0000;
		notes[72] = 4'b0001;  //measure 18
		notes[73] = 4'b0010;
		notes[74] = 4'b1000;
		notes[75] = 4'b0001;  
		notes[76] = 4'b1000;  //measure 19
		notes[77] = 4'b0010;
		notes[78] = 4'b0001;
		notes[79] = 4'b1000;
		notes[80] = 4'b0001;  //measure 20
		notes[81] = 4'b0010;
		notes[82] = 4'b1000;
		notes[83] = 4'b0001;
		notes[84] = 4'b0100;  //measure 21
		notes[85] = 4'b0010;
		notes[86] = 4'b0001;
		notes[87] = 4'b1000;
		notes[88] = 4'b0001;  //measure 22
		notes[89] = 4'b0100;
		notes[90] = 4'b0010;
		notes[91] = 4'b0000;
		notes[92] = 4'b0000;  //measure 23
		notes[93] = 4'b0010;
		notes[94] = 4'b0001;
		notes[95] = 4'b1000;
		notes[96] = 4'b0010;  //measure 24
		notes[97] = 4'b0100;
		notes[98] = 4'b0010;
		notes[99] = 4'b1000;
		notes[100] = 4'b0001;  //measure 25
		notes[101] = 4'b0001;
		notes[102] = 4'b1000;
		notes[103] = 4'b0001;
		notes[104] = 4'b0100;  //measure 26
		notes[105] = 4'b0010;
		notes[106] = 4'b1000;
		notes[107] = 4'b0001;
		notes[108] = 4'b0100;  //measure 27
		notes[109] = 4'b0100;
		notes[110] = 4'b1000;
		notes[111] = 4'b0100;
		notes[112] = 4'b0001;  //measure 28
		notes[113] = 4'b1000;
		notes[114] = 4'b0010;
		notes[115] = 4'b0001; 
		notes[116] = 4'b0001;  //measure 29
		notes[117] = 4'b1000;
		notes[118] = 4'b1000;
		notes[119] = 4'b0010;
		notes[120] = 4'b1000;  //measure 30
		notes[121] = 4'b0001;
		notes[122] = 4'b1001;
		notes[123] = 4'b1100;
		notes[124] = 4'b0100;  //measure 31
		notes[125] = 4'b1000;
		notes[126] = 4'b1000;
		notes[127] = 4'b0100;
		notes[128] = 4'b0100;  //measure 32
		notes[129] = 4'b1000;
		notes[130] = 4'b0010;
		notes[131] = 4'b0100;
		notes[132] = 4'b0100;  //measure 33
		notes[133] = 4'b0001;
		notes[134] = 4'b0001;
		notes[135] = 4'b0100;
		notes[136] = 4'b0100;  //measure 34
		notes[137] = 4'b0001;
		notes[138] = 4'b0100;
		notes[139] = 4'b0001;
		notes[140] = 4'b0000;  //measure 35
		notes[141] = 4'b0001;
		notes[142] = 4'b0000;
		notes[143] = 4'b0000;
		notes[144] = 4'b0000;  //measure 36
		notes[145] = 4'b0000;
		notes[146] = 4'b0000;
		notes[147] = 4'b0000;
		notes[148] = 4'b0000;  //measure 37
		notes[149] = 4'b0010;
		notes[150] = 4'b0100;
		notes[151] = 4'b0001;
		notes[152] = 4'b0000;  //measure 38
		notes[153] = 4'b0000;
		notes[154] = 4'b0001;
		notes[155] = 4'b0100;
		notes[156] = 4'b1000;  //measure 39
		notes[157] = 4'b0001;
		notes[158] = 4'b0001;
		notes[159] = 4'b0100;
		notes[160] = 4'b0000;  //measure 40
		notes[161] = 4'b0000;
		notes[162] = 4'b0100;
		notes[163] = 4'b0001;
		notes[164] = 4'b1000;  //measure 41
		notes[165] = 4'b0001;
		notes[166] = 4'b0001;
		notes[167] = 4'b0010;
		notes[168] = 4'b1000;  //measure 42
		notes[169] = 4'b0010;
		notes[170] = 4'b0001;
		notes[171] = 4'b1000;
		notes[172] = 4'b0010;  //measure 43
		notes[173] = 4'b0100;
		notes[174] = 4'b0100;
		notes[175] = 4'b0001;
		notes[176] = 4'b0100;  //measure 44
		notes[177] = 4'b0010;
		notes[178] = 4'b1000;
		notes[179] = 4'b0010;
		notes[180] = 4'b0001;  //measure 45
		notes[181] = 4'b1000;
		notes[182] = 4'b1000;
		notes[183] = 4'b0001;  
		notes[184] = 4'b0000;  //measure 46
		notes[185] = 4'b0000;
		notes[186] = 4'b0001;
		notes[187] = 4'b0100;
		notes[188] = 4'b0001;  //measure 47
		notes[189] = 4'b1000;
		notes[190] = 4'b1000;
		notes[191] = 4'b0010;
		notes[192] = 4'b0000;  //measure 48
		notes[193] = 4'b0000;
		notes[194] = 4'b0010;
		notes[195] = 4'b0001;
		notes[196] = 4'b1000;  //measure 49
		notes[197] = 4'b0100;
		notes[198] = 4'b0100;
		notes[199] = 4'b0001;				
		notes[200] = 4'b0100;  //measure 50
		notes[201] = 4'b0100;
		notes[202] = 4'b0000;
		notes[203] = 4'b1000;
		notes[204] = 4'b0010;  //measure 51
		notes[205] = 4'b0001;
		notes[206] = 4'b0001;
		notes[207] = 4'b1000;
		notes[208] = 4'b1001;  //measure 52
		notes[209] = 4'b0101;
		notes[210] = 4'b0100;
		notes[211] = 4'b0000;
		notes[212] = 4'b0000;  //measure 53
		notes[213] = 4'b0010;
		notes[214] = 4'b1000;
		notes[215] = 4'b0100;
		notes[216] = 4'b0001;  //measure 54
		notes[217] = 4'b0010;
		notes[218] = 4'b1000;
		notes[219] = 4'b0100;
		notes[220] = 4'b0100;  //measure 55
		notes[221] = 4'b1000;
		notes[222] = 4'b0001;
		notes[223] = 4'b0010;
		notes[224] = 4'b1000;  //measure 56
		notes[225] = 4'b0100;
		notes[226] = 4'b0000;
		notes[227] = 4'b0000;
		notes[228] = 4'b0000;  //measure 57
		notes[229] = 4'b0000;
		notes[230] = 4'b0100;
		notes[231] = 4'b0001;  //last beat of last measure
		notes[232] = 4'b0000;  //measure 58 
		notes[233] = 4'b0000;
		notes[234] = 4'b0000;
		notes[235] = 4'b0000;
		notes[236] = 4'b0000;  //measure 59
		notes[237] = 4'b0000;
		notes[238] = 4'b0000;
		notes[239] = 4'b0000;
		notes[240] = 4'b0000;  //measure 60
		notes[241] = 4'b0000;
		notes[242] = 4'b0000;
		notes[243] = 4'b0000;
		notes[244] = 4'b0000;  //measure 61
		notes[245] = 4'b0000;
		notes[246] = 4'b0000;
		notes[247] = 4'b0000;
		notes[248] = 4'b0000;  //measure 62
		notes[249] = 4'b0000;
		notes[250] = 4'b0000;
		notes[251] = 4'b0000;
		notes[252] = 4'b0000;  //measure 63
		notes[253] = 4'b0000;
		notes[254] = 4'b0000;
		notes[255] = 4'b0000;
	
end

always @(posedge clk) begin
		data = notes[addr];
end

endmodule